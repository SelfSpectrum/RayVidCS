CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
9 2-In AND~
219 249 597 0 3 22
0 4 5 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7876 0 0
2
5.90075e-315 0
0
14 Logic Display~
6 1028 46 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.90075e-315 0
0
8 2-In OR~
219 360 544 0 3 22
0 7 5 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9172 0 0
2
5.90075e-315 0
0
5 7415~
219 248 527 0 4 22
0 4 8 9 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 5 0
1 U
7100 0 0
2
5.90075e-315 0
0
8 2-In OR~
219 242 266 0 3 22
0 9 5 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3820 0 0
2
5.90075e-315 0
0
8 2-In OR~
219 358 488 0 3 22
0 11 5 12
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7678 0 0
2
5.90075e-315 0
0
8 2-In OR~
219 525 414 0 3 22
0 14 12 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
961 0 0
2
5.90075e-315 0
0
14 Logic Display~
6 992 48 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
45051.5 0
0
14 Logic Display~
6 954 49 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
45051.5 1
0
14 Logic Display~
6 908 51 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
45051.5 2
0
14 Logic Display~
6 864 53 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
45051.5 3
0
14 Logic Display~
6 817 54 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
45051.5 4
0
14 Logic Display~
6 765 53 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
45051.5 5
0
14 Logic Display~
6 707 55 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
45051.5 6
0
8 2-In OR~
219 387 275 0 3 22
0 10 2 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9424 0 0
2
45051.5 7
0
8 2-In OR~
219 517 97 0 3 22
0 4 16 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9968 0 0
2
45051.5 8
0
14 Logic Display~
6 627 57 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
45051.5 9
0
8 2-In OR~
219 380 154 0 3 22
0 8 10 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8464 0 0
2
45051.5 10
0
9 2-In AND~
219 246 461 0 3 22
0 9 8 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7168 0 0
2
45051.5 11
0
9 2-In AND~
219 248 403 0 3 22
0 9 4 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3171 0 0
2
45051.5 12
0
9 2-In AND~
219 250 340 0 3 22
0 4 8 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4139 0 0
2
45051.5 13
0
8 Hex Key~
166 148 103 0 11 12
0 4 8 9 5 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6435 0 0
2
45051.5 14
0
34
3 2 2 0 0 4224 0 21 15 0 0 4
271 340
366 340
366 284
374 284
3 1 3 0 0 4224 0 1 2 0 0 3
270 597
1028 597
1028 64
1 1 4 0 0 8320 0 1 22 0 0 3
225 588
157 588
157 127
4 2 5 0 0 4096 0 22 1 0 0 3
139 127
139 606
225 606
3 1 6 0 0 4224 0 3 9 0 0 3
393 544
954 544
954 67
4 1 7 0 0 4224 0 4 3 0 0 4
269 527
339 527
339 535
347 535
4 2 5 0 0 0 0 22 3 0 0 3
139 127
139 553
347 553
1 1 4 0 0 0 0 22 4 0 0 3
157 127
157 518
224 518
2 2 8 0 0 4224 0 22 4 0 0 3
151 127
151 527
224 527
3 3 9 0 0 4224 0 22 4 0 0 3
145 127
145 536
224 536
1 4 5 0 0 8320 0 8 22 0 0 4
992 66
992 192
139 192
139 127
3 1 10 0 0 12416 0 5 12 0 0 5
275 266
360 266
360 212
817 212
817 72
3 2 10 0 0 0 0 5 18 0 0 4
275 266
360 266
360 163
367 163
3 1 10 0 0 0 0 5 15 0 0 2
275 266
374 266
3 1 9 0 0 0 0 22 5 0 0 3
145 127
145 257
229 257
4 2 5 0 0 0 0 22 5 0 0 3
139 127
139 275
229 275
4 2 5 0 0 0 0 22 6 0 0 3
139 127
139 497
345 497
3 1 11 0 0 4224 0 19 6 0 0 4
267 461
337 461
337 479
345 479
3 1 12 0 0 4224 0 6 10 0 0 3
391 488
908 488
908 69
3 2 12 0 0 0 0 6 7 0 0 4
391 488
504 488
504 423
512 423
3 1 13 0 0 8320 0 7 11 0 0 3
558 414
864 414
864 71
3 1 14 0 0 4224 0 20 7 0 0 4
269 403
496 403
496 405
512 405
3 1 15 0 0 4224 0 15 13 0 0 3
420 275
765 275
765 71
3 1 16 0 0 4224 0 18 14 0 0 3
413 154
707 154
707 73
3 1 17 0 0 4224 0 16 17 0 0 3
550 97
627 97
627 75
3 2 16 0 0 0 0 18 16 0 0 4
413 154
496 154
496 106
504 106
1 1 4 0 0 0 0 22 16 0 0 5
157 127
157 131
364 131
364 88
504 88
2 1 8 0 0 0 0 22 18 0 0 3
151 127
151 145
367 145
2 2 8 0 0 0 0 19 22 0 0 3
222 470
151 470
151 127
3 1 9 0 0 0 0 22 19 0 0 3
145 127
145 452
222 452
2 1 4 0 0 0 0 20 22 0 0 3
224 412
157 412
157 127
3 1 9 0 0 0 0 22 20 0 0 3
145 127
145 394
224 394
2 2 8 0 0 0 0 22 21 0 0 3
151 127
151 349
226 349
1 1 4 0 0 0 0 22 21 0 0 3
157 127
157 331
226 331
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
376 259 413 283
386 267 402 283
2 L3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
506 82 543 106
516 90 532 106
2 L1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
369 138 406 162
379 146 395 162
2 L2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
226 447 263 471
236 455 252 471
2 BC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
229 388 266 412
239 396 255 412
2 BD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
228 323 265 347
238 331 254 347
2 CD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
515 396 552 420
525 404 541 420
2 L5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
346 471 383 495
356 479 372 495
2 L6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
231 250 268 274
241 258 257 274
2 L4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
222 511 267 535
232 519 256 535
3 BCD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
349 528 386 552
359 536 375 552
2 L7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
229 582 266 606
239 590 255 606
2 L9
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
