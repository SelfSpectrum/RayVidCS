CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
140 120 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 394 1364 707
42991634 0
0
6 Title:
5 Name:
0
0
0
14
9 2-In AND~
219 568 568 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
5130 0 0
2
45072.8 0
0
9 2-In AND~
219 568 475 0 3 22
0 9 8 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
391 0 0
2
45072.8 0
0
9 2-In AND~
219 567 395 0 3 22
0 7 6 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3124 0 0
2
45072.7 0
0
8 2-In OR~
219 551 279 0 3 22
0 11 10 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3421 0 0
2
45072.7 0
0
14 Logic Display~
6 1107 94 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-6 -21 8 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
8157 0 0
2
45072.7 0
0
14 Logic Display~
6 1014 96 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
5572 0 0
2
45072.7 0
0
14 Logic Display~
6 989 87 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
8901 0 0
2
45072.7 0
0
14 Logic Display~
6 839 39 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
45072.7 0
0
14 Logic Display~
6 796 39 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
4747 0 0
2
45072.7 0
0
14 Logic Display~
6 748 32 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
45072.7 0
0
14 Logic Display~
6 666 45 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
45072.7 0
0
4 4028
219 168 457 0 14 29
0 12 13 14 15 10 6 8 20 21
22 23 24 25 26
0
0 0 4848 0
4 4028
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 10 3 14 2 15 1
6 7 4 9 5 11 12 13 10 3
14 2 15 1 6 7 4 9 5 0
65 0 0 512 0 0 0 0
1 U
9998 0 0
2
45072.7 0
0
4 4028
219 164 225 0 14 29
0 12 13 14 15 11 7 9 27 28
29 30 31 32 33
0
0 0 4848 0
4 4028
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 10 3 14 2 15 1
6 7 4 9 5 11 12 13 10 3
14 2 15 1 6 7 4 9 5 0
65 0 0 512 0 0 0 0
1 U
3536 0 0
2
45072.7 0
0
8 Hex Key~
166 56 165 0 11 12
0 15 14 13 12 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
4597 0 0
2
45072.7 0
0
21
3 1 0 0 0 0 0 1 5 0 0 3
589 568
1107 568
1107 112
3 1 0 0 0 0 0 1 11 0 0 3
589 568
666 568
666 63
1 8 0 0 0 16 0 1 13 0 0 4
544 559
443 559
443 243
196 243
8 2 0 0 0 0 0 12 1 0 0 4
200 475
310 475
310 577
544 577
1 3 0 0 0 0 0 8 2 0 0 3
839 57
839 475
589 475
7 2 8 0 0 12416 0 12 2 0 0 2
200 484
544 484
7 1 9 0 0 8320 0 13 2 0 0 4
196 252
393 252
393 466
544 466
3 1 2 0 0 128 0 3 10 0 0 3
588 395
748 395
748 50
6 2 6 0 0 12416 0 12 3 0 0 4
200 493
268 493
268 404
543 404
6 1 7 0 0 128 0 13 3 0 0 4
196 261
426 261
426 386
543 386
1 3 5 0 0 128 0 11 4 0 0 3
666 63
666 279
584 279
5 2 10 0 0 12416 0 12 4 0 0 4
200 502
235 502
235 288
538 288
5 1 11 0 0 4224 0 13 4 0 0 2
196 270
538 270
1 4 12 0 0 8320 0 12 14 0 0 3
136 475
47 475
47 189
3 2 13 0 0 4224 0 14 12 0 0 3
53 189
53 484
136 484
3 2 14 0 0 8320 0 12 14 0 0 3
136 493
59 493
59 189
1 4 15 0 0 4224 0 14 12 0 0 3
65 189
65 502
136 502
1 4 12 0 0 128 0 13 14 0 0 3
132 243
47 243
47 189
2 3 13 0 0 128 0 13 14 0 0 3
132 252
53 252
53 189
3 2 14 0 0 128 0 13 14 0 0 3
132 261
59 261
59 189
1 4 15 0 0 128 0 14 13 0 0 3
65 189
65 270
132 270
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
543 553 588 577
553 561 577 577
3 A-B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
543 460 588 484
553 468 577 484
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
535 381 596 405
545 389 585 405
5 AandB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
533 263 586 287
543 271 575 287
4 AorB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1066 42 1151 66
1076 50 1140 66
8 overflow
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
