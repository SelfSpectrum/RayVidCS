CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 540 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 60 695 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3951 0 0
2
5.90079e-315 0
0
13 Logic Switch~
5 60 567 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8885 0 0
2
5.90079e-315 0
0
13 Logic Switch~
5 792 63 0 1 11
0 30
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
5.90079e-315 0
0
9 Inverter~
13 210 683 0 2 22
0 5 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
9265 0 0
2
5.90079e-315 0
0
9 Inverter~
13 195 760 0 2 22
0 4 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
9442 0 0
2
5.90079e-315 0
0
9 Inverter~
13 192 719 0 2 22
0 2 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
9424 0 0
2
5.90079e-315 0
0
9 Inverter~
13 190 661 0 2 22
0 6 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9968 0 0
2
5.90079e-315 0
0
12 Hex Display~
7 1108 100 0 18 19
10 39 38 37 36 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9281 0 0
2
5.90079e-315 0
0
12 Hex Display~
7 1041 103 0 16 19
10 26 25 24 23 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8464 0 0
2
5.90079e-315 0
0
8 Hex Key~
166 201 29 0 11 12
0 27 28 29 48 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
7168 0 0
2
5.90079e-315 0
0
8 Hex Key~
166 146 56 0 11 12
0 6 5 2 4 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3171 0 0
2
5.90079e-315 0
0
8 Hex Key~
166 87 58 0 11 12
0 9 8 3 7 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4139 0 0
2
5.90079e-315 0
0
7 74LS251
144 714 551 0 14 29
0 10 8 4 10 10 31 10 10 29
28 27 30 49 26
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U13
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6435 0 0
2
5.90079e-315 0
0
7 74LS251
144 713 448 0 14 29
0 10 9 2 10 18 32 40 44 29
28 27 30 50 36
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U12
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5283 0 0
2
5.90079e-315 0
0
7 74LS251
144 717 765 0 14 29
0 10 7 8 10 10 10 10 10 29
28 27 30 51 24
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6874 0 0
2
5.90079e-315 0
0
7 74LS251
144 704 150 0 14 29
0 10 5 10 13 21 35 43 47 29
28 27 30 52 39
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
3 U10
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
5305 0 0
2
5.90079e-315 0
0
7 74LS251
144 717 664 0 14 29
0 10 3 9 10 10 10 10 10 29
28 27 30 53 25
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.90079e-315 0
0
7 74LS251
144 717 872 0 14 29
0 10 10 3 10 10 10 10 10 29
28 27 30 54 23
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
969 0 0
2
5.90079e-315 0
0
7 74LS251
144 710 341 0 14 29
0 10 4 5 11 19 33 41 45 29
28 27 30 55 37
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8402 0 0
2
5.90079e-315 0
0
4 4008
219 337 661 0 14 29
0 7 3 8 9 14 15 16 17 22
21 20 19 18 56
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U7
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3751 0 0
2
5.90079e-315 0
0
4 4008
219 337 527 0 14 29
0 7 3 8 9 4 2 5 6 10
35 34 33 32 31
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U6
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 1 0 0 0
1 U
4292 0 0
2
5.90079e-315 0
0
7 74LS251
144 707 246 0 14 29
0 10 2 6 12 20 34 42 46 29
28 27 30 57 38
0
0 0 4848 0
7 74LS251
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 9
10 11 7 6 5 12 13 14 15 1
2 3 4 9 10 11 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6118 0 0
2
5.90079e-315 0
0
6 74LS85
106 336 805 0 14 29
0 7 3 8 9 4 2 5 6 58
59 60 11 12 13
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
34 0 0
2
5.90079e-315 0
0
9 2-In AND~
219 341 424 0 3 22
0 6 9 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6357 0 0
2
5.90079e-315 0
0
9 2-In AND~
219 339 382 0 3 22
0 5 8 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
319 0 0
2
5.90079e-315 0
0
9 2-In AND~
219 341 338 0 3 22
0 2 3 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3976 0 0
2
5.90079e-315 0
0
9 2-In AND~
219 342 296 0 3 22
0 4 7 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7634 0 0
2
5.90079e-315 0
0
8 2-In OR~
219 332 229 0 3 22
0 6 9 47
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
523 0 0
2
5.90079e-315 0
0
8 2-In OR~
219 333 187 0 3 22
0 5 8 46
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6748 0 0
2
5.90079e-315 0
0
8 2-In OR~
219 332 148 0 3 22
0 2 3 45
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6901 0 0
2
5.90079e-315 0
0
8 2-In OR~
219 332 107 0 3 22
0 4 7 44
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
842 0 0
2
5.90079e-315 0
0
150
2 5 0 0 0 0 0 7 20 0 0 2
211 661
305 661
2 6 0 0 0 0 0 4 20 0 0 4
231 683
234 683
234 670
305 670
2 7 0 0 0 0 0 6 20 0 0 4
213 719
243 719
243 679
305 679
2 8 0 0 0 0 0 5 20 0 0 4
216 760
255 760
255 688
305 688
1 0 0 0 0 0 0 5 0 0 62 4
180 760
160 760
160 761
155 761
0 1 0 0 0 0 0 0 6 61 0 2
149 719
177 719
0 1 0 0 0 0 0 0 4 60 0 2
143 683
195 683
0 1 0 0 0 0 0 0 7 59 0 2
137 661
175 661
1 3 2 0 0 4096 0 30 11 0 0 3
319 139
143 139
143 80
2 3 3 0 0 4096 0 30 12 0 0 3
319 157
84 157
84 82
4 1 4 0 0 4096 0 11 27 0 0 3
137 80
137 287
318 287
1 3 2 0 0 8192 0 26 11 0 0 3
317 329
143 329
143 80
1 2 5 0 0 8192 0 25 11 0 0 3
315 373
149 373
149 80
1 1 6 0 0 4096 0 11 24 0 0 3
155 80
155 415
317 415
4 2 7 0 0 8192 0 12 27 0 0 3
78 82
78 305
318 305
3 2 3 0 0 4096 0 12 26 0 0 3
84 82
84 347
317 347
2 2 8 0 0 4096 0 12 25 0 0 3
90 82
90 391
315 391
2 1 9 0 0 8192 0 24 12 0 0 3
317 433
96 433
96 82
1 2 10 0 0 4096 0 18 18 0 0 2
685 845
685 854
1 2 7 0 0 12288 0 21 15 0 0 4
305 491
271 491
271 747
685 747
2 2 3 0 0 12288 0 21 17 0 0 6
305 500
276 500
276 712
662 712
662 646
685 646
3 2 8 0 0 12288 0 21 13 0 0 6
305 509
291 509
291 593
664 593
664 533
682 533
2 4 9 0 0 0 0 14 21 0 0 6
681 430
373 430
373 471
297 471
297 518
305 518
4 2 4 0 0 8192 0 11 19 0 0 5
137 80
137 318
660 318
660 323
678 323
3 2 2 0 0 8192 0 11 22 0 0 5
143 80
143 209
667 209
667 228
675 228
2 2 5 0 0 8192 0 11 16 0 0 5
149 80
149 128
654 128
654 132
672 132
1 3 10 0 0 8192 0 16 16 0 0 4
672 123
664 123
664 141
672 141
2 3 3 0 0 12288 0 23 18 0 0 4
304 787
290 787
290 863
685 863
3 3 8 0 0 12288 0 23 15 0 0 4
304 796
295 796
295 756
685 756
4 3 9 0 0 12304 0 23 17 0 0 6
304 805
301 805
301 723
637 723
637 655
685 655
4 1 10 0 0 8192 0 14 14 0 0 4
681 448
658 448
658 421
681 421
4 3 4 0 0 8192 0 11 13 0 0 5
137 80
137 583
669 583
669 542
682 542
3 3 2 0 0 8192 0 11 14 0 0 5
143 80
143 444
673 444
673 439
681 439
2 3 5 0 0 8192 0 11 19 0 0 5
149 80
149 318
670 318
670 332
678 332
1 3 6 0 0 8192 0 11 22 0 0 5
155 80
155 249
667 249
667 237
675 237
1 1 10 0 0 8192 0 22 16 0 0 4
675 219
659 219
659 123
672 123
1 1 10 0 0 0 0 19 22 0 0 4
678 314
662 314
662 219
675 219
1 1 10 0 0 8192 0 14 19 0 0 4
681 421
665 421
665 314
678 314
1 1 10 0 0 0 0 13 14 0 0 4
682 524
668 524
668 421
681 421
4 1 10 0 0 0 0 13 13 0 0 4
682 551
674 551
674 524
682 524
4 1 10 0 0 0 0 17 17 0 0 4
685 664
672 664
672 637
685 637
4 1 10 0 0 0 0 15 15 0 0 4
685 765
658 765
658 738
685 738
4 1 10 0 0 0 0 18 18 0 0 4
685 872
672 872
672 845
685 845
4 5 10 0 0 0 0 17 17 0 0 2
685 664
685 673
5 4 10 0 0 0 0 18 18 0 0 2
685 881
685 872
5 4 10 0 0 0 0 15 15 0 0 2
685 774
685 765
5 4 10 0 0 0 0 13 13 0 0 2
682 560
682 551
12 4 11 0 0 8320 0 23 19 0 0 4
368 823
510 823
510 341
678 341
13 4 12 0 0 8320 0 23 22 0 0 4
368 832
502 832
502 246
675 246
14 4 13 0 0 8320 0 23 16 0 0 4
368 841
497 841
497 150
672 150
6 5 10 0 0 0 0 18 18 0 0 2
685 890
685 881
6 5 10 0 0 0 0 15 15 0 0 2
685 783
685 774
6 5 10 0 0 0 0 17 17 0 0 2
685 682
685 673
7 5 10 0 0 0 0 13 13 0 0 4
682 578
623 578
623 560
682 560
13 5 18 0 0 12416 0 20 14 0 0 4
369 643
489 643
489 457
681 457
12 5 19 0 0 8320 0 20 19 0 0 4
369 652
481 652
481 350
678 350
11 5 20 0 0 8320 0 20 22 0 0 4
369 661
468 661
468 255
675 255
10 5 21 0 0 8320 0 20 16 0 0 4
369 670
460 670
460 159
672 159
4 5 4 0 0 4224 0 11 23 0 0 3
137 80
137 814
304 814
6 3 2 0 0 8320 0 23 11 0 0 3
304 823
143 823
143 80
2 7 5 0 0 4224 0 11 23 0 0 3
149 80
149 832
304 832
8 1 6 0 0 8320 0 23 11 0 0 3
304 841
155 841
155 80
1 4 9 0 0 4224 0 12 23 0 0 3
96 82
96 805
304 805
3 2 8 0 0 8320 0 23 12 0 0 3
304 796
90 796
90 82
3 2 3 0 0 4224 0 12 23 0 0 3
84 82
84 787
304 787
1 4 7 0 0 8320 0 23 12 0 0 3
304 778
78 778
78 82
4 1 7 0 0 0 0 12 20 0 0 3
78 82
78 625
305 625
2 3 3 0 0 0 0 20 12 0 0 3
305 634
84 634
84 82
2 3 8 0 0 0 0 12 20 0 0 3
90 82
90 643
305 643
4 1 9 0 0 0 0 20 12 0 0 3
305 652
96 652
96 82
1 9 22 0 0 8320 0 1 20 0 0 3
72 695
72 697
305 697
7 6 10 0 0 0 0 18 18 0 0 2
685 899
685 890
7 6 10 0 0 0 0 15 15 0 0 2
685 792
685 783
7 6 10 0 0 0 0 17 17 0 0 2
685 691
685 682
8 7 10 0 0 0 0 18 18 0 0 2
685 908
685 899
8 8 10 0 0 0 0 15 18 0 0 4
685 801
677 801
677 908
685 908
8 7 10 0 0 0 0 15 15 0 0 2
685 801
685 792
8 8 10 0 0 0 0 17 15 0 0 4
685 700
672 700
672 801
685 801
8 7 10 0 0 0 0 17 17 0 0 2
685 700
685 691
8 7 10 0 0 0 0 13 13 0 0 2
682 587
682 578
8 8 10 0 0 8192 0 13 17 0 0 4
682 587
677 587
677 700
685 700
1 8 10 0 0 12416 0 2 13 0 0 4
72 567
301 567
301 587
682 587
14 4 23 0 0 8320 0 18 9 0 0 3
749 908
1032 908
1032 127
14 3 24 0 0 8320 0 15 9 0 0 3
749 801
1038 801
1038 127
14 2 25 0 0 8320 0 17 9 0 0 3
749 700
1044 700
1044 127
14 1 26 0 0 8320 0 13 9 0 0 3
746 587
1050 587
1050 127
11 11 27 0 0 8192 0 15 18 0 0 4
749 756
788 756
788 863
749 863
10 10 28 0 0 8192 0 18 15 0 0 4
749 854
783 854
783 747
749 747
9 9 29 0 0 8192 0 15 18 0 0 4
749 738
773 738
773 845
749 845
9 9 29 0 0 0 0 17 15 0 0 4
749 637
793 637
793 738
749 738
10 10 28 0 0 0 0 15 17 0 0 4
749 747
788 747
788 646
749 646
11 11 27 0 0 0 0 17 15 0 0 4
749 655
778 655
778 756
749 756
9 9 29 0 0 8192 0 13 17 0 0 4
746 524
788 524
788 637
749 637
10 10 28 0 0 8192 0 13 17 0 0 4
746 533
783 533
783 646
749 646
11 11 27 0 0 8192 0 13 17 0 0 4
746 542
773 542
773 655
749 655
12 12 30 0 0 8192 0 15 18 0 0 4
755 765
768 765
768 872
755 872
12 12 30 0 0 0 0 17 15 0 0 4
755 664
763 664
763 765
755 765
12 12 30 0 0 8320 0 13 17 0 0 4
752 551
768 551
768 664
755 664
12 12 30 0 0 0 0 14 13 0 0 4
751 448
765 448
765 551
752 551
9 9 29 0 0 0 0 14 13 0 0 4
745 421
785 421
785 524
746 524
10 10 28 0 0 0 0 14 13 0 0 4
745 430
780 430
780 533
746 533
11 11 27 0 0 0 0 14 13 0 0 4
745 439
760 439
760 542
746 542
14 6 31 0 0 4224 0 21 13 0 0 4
369 491
644 491
644 569
682 569
13 6 32 0 0 12416 0 21 14 0 0 4
369 509
453 509
453 466
681 466
12 6 33 0 0 12416 0 21 19 0 0 4
369 518
448 518
448 359
678 359
11 6 34 0 0 8320 0 21 22 0 0 4
369 527
440 527
440 264
675 264
10 6 35 0 0 8320 0 21 16 0 0 4
369 536
431 536
431 168
672 168
1 9 10 0 0 0 0 2 21 0 0 4
72 567
297 567
297 563
305 563
1 4 7 0 0 0 0 21 12 0 0 3
305 491
78 491
78 82
2 3 3 0 0 0 0 21 12 0 0 3
305 500
84 500
84 82
3 2 8 0 0 0 0 21 12 0 0 3
305 509
90 509
90 82
4 1 9 0 0 0 0 21 12 0 0 3
305 518
96 518
96 82
5 4 4 0 0 0 0 21 11 0 0 3
305 527
137 527
137 80
6 3 2 0 0 0 0 21 11 0 0 3
305 536
143 536
143 80
2 7 5 0 0 0 0 11 21 0 0 3
149 80
149 545
305 545
1 8 6 0 0 0 0 11 21 0 0 3
155 80
155 554
305 554
14 4 36 0 0 4224 0 14 8 0 0 3
745 484
1099 484
1099 124
14 3 37 0 0 4224 0 19 8 0 0 3
742 377
1105 377
1105 124
14 2 38 0 0 4224 0 22 8 0 0 3
739 282
1111 282
1111 124
14 1 39 0 0 4224 0 16 8 0 0 5
736 186
984 186
984 185
1117 185
1117 124
9 9 29 0 0 0 0 14 19 0 0 4
745 421
782 421
782 314
742 314
10 10 28 0 0 0 0 14 19 0 0 4
745 430
767 430
767 323
742 323
11 11 27 0 0 0 0 19 14 0 0 4
742 332
776 332
776 439
745 439
9 9 29 0 0 0 0 22 19 0 0 4
739 219
787 219
787 314
742 314
10 10 28 0 0 0 0 19 22 0 0 4
742 323
776 323
776 228
739 228
11 11 27 0 0 0 0 22 19 0 0 4
739 237
762 237
762 332
742 332
12 12 30 0 0 0 0 19 14 0 0 4
748 341
771 341
771 448
751 448
12 12 30 0 0 0 0 22 19 0 0 4
745 246
757 246
757 341
748 341
12 12 30 0 0 0 0 16 22 0 0 4
742 150
781 150
781 246
745 246
1 12 30 0 0 0 0 3 16 0 0 3
792 75
792 150
742 150
9 9 29 0 0 0 0 16 22 0 0 4
736 123
776 123
776 219
739 219
10 10 28 0 0 0 0 16 22 0 0 4
736 132
771 132
771 228
739 228
11 11 27 0 0 0 0 16 22 0 0 4
736 141
766 141
766 237
739 237
3 7 40 0 0 12416 0 27 14 0 0 4
363 296
402 296
402 475
681 475
3 7 41 0 0 12416 0 26 19 0 0 4
362 338
407 338
407 368
678 368
3 7 42 0 0 12416 0 25 22 0 0 4
360 382
412 382
412 273
675 273
3 7 43 0 0 12416 0 24 16 0 0 4
362 424
419 424
419 177
672 177
3 9 29 0 0 8320 0 10 16 0 0 5
198 53
198 79
760 79
760 123
736 123
2 10 28 0 0 8320 0 10 16 0 0 5
204 53
204 70
755 70
755 132
736 132
1 11 27 0 0 8320 0 10 16 0 0 5
210 53
210 61
750 61
750 141
736 141
3 8 44 0 0 8320 0 31 14 0 0 4
365 107
392 107
392 484
681 484
3 8 45 0 0 12416 0 30 19 0 0 4
365 148
388 148
388 377
678 377
3 8 46 0 0 12416 0 29 22 0 0 4
366 187
381 187
381 282
675 282
3 8 47 0 0 12416 0 28 16 0 0 5
365 229
376 229
376 194
672 194
672 186
4 2 7 0 0 0 0 12 31 0 0 3
78 82
78 116
319 116
4 1 4 0 0 0 0 11 31 0 0 3
137 80
137 98
319 98
2 2 8 0 0 0 0 12 29 0 0 5
90 82
90 194
307 194
307 196
320 196
2 1 5 0 0 0 0 11 29 0 0 3
149 80
149 178
320 178
1 1 6 0 0 0 0 11 28 0 0 3
155 80
155 220
319 220
1 2 9 0 0 0 0 12 28 0 0 5
96 82
96 237
311 237
311 238
319 238
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
73 -4 102 20
83 4 91 20
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
131 -6 160 18
141 2 149 18
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
218 6 247 30
228 14 236 30
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
314 42 357 57
328 53 342 64
2 Or
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
314 243 364 258
328 254 349 265
3 and
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
306 444 356 459
320 456 341 467
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
310 573 360 588
324 584 345 595
3 A-B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
310 711 360 726
324 723 345 734
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1168 121 1269 145
1179 130 1257 146
13 1 A mayor a B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1177 95 1266 119
1188 104 1254 120
11 2 A igual B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1173 72 1274 96
1184 80 1262 96
13 4 B mayor a A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
